type memoryPicture is array(0 to 14, 0 to 14) of integer;
constant picture : memoryPicture:=(
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#20#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#c3#,16#c3#,16#0#,16#0#,16#c3#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#c3#,16#c3#,16#c3#,16#0#,16#c3#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#20#,16#0#,16#c3#,16#c3#,16#0#,16#c3#,16#c3#,16#0#,16#c3#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#c3#,16#c3#,16#c3#,16#c3#,16#c3#,16#0#,16#c3#,16#20#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#c3#,16#c3#,16#c3#,16#c3#,16#c3#,16#0#,16#c3#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#c3#,16#c3#,16#c3#,16#c3#,16#c3#,16#0#,16#c3#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#c3#,16#c3#,16#0#,16#c3#,16#c3#,16#0#,16#c3#,16#4#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#c3#,16#c3#,16#c3#,16#0#,16#c3#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#c3#,16#c3#,16#0#,16#0#,16#c3#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#20#,16#0#),
(16#0#,16#0#,16#4#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#));