type memoryPicture is array(0 to 199, 0 to 149) of integer;
constant picture : memoryPicture:=(
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#0#,16#4#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#4#,16#fb#,16#20#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#1#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#4#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#20#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#20#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#d7#,16#d7#,16#d7#,16#d7#,16#d7#,16#d7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#ff#,16#ff#,16#0#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#20#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#0#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#20#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#ff#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#18#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#0#,16#ff#,16#ff#,16#bb#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#14#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#9b#,16#ff#,16#0#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#0#,16#18#,16#18#,16#14#,16#18#,16#18#,16#14#,16#14#,16#18#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#9b#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#0#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#ff#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#b8#,16#bc#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#d7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#20#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#b8#,16#bc#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#0#,16#18#,16#bc#,16#b8#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#0#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#14#,16#18#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#0#,16#18#,16#18#,16#14#,16#18#,16#18#,16#18#,16#18#,16#18#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#d7#,16#b7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#18#,16#14#,16#18#,16#14#,16#18#,16#18#,16#18#,16#18#,16#0#,16#18#,16#18#,16#14#,16#14#,16#14#,16#14#,16#18#,16#18#,16#18#,16#18#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#4#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#ff#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#18#,16#18#,16#18#,16#18#,16#18#,16#14#,16#18#,16#14#,16#0#,16#14#,16#18#,16#14#,16#18#,16#18#,16#14#,16#18#,16#14#,16#14#,16#18#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#0#,16#ff#,16#ff#,16#bb#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#18#,16#14#,16#18#,16#18#,16#18#,16#18#,16#14#,16#18#,16#0#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#18#,16#18#,16#18#,16#18#,16#14#,16#18#,16#14#,16#14#,16#0#,16#18#,16#14#,16#18#,16#18#,16#18#,16#18#,16#14#,16#18#,16#18#,16#18#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#20#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#18#,16#18#,16#14#,16#18#,16#18#,16#18#,16#18#,16#18#,16#0#,16#14#,16#14#,16#14#,16#18#,16#18#,16#14#,16#14#,16#14#,16#18#,16#18#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#ff#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#18#,16#18#,16#18#,16#18#,16#14#,16#18#,16#14#,16#38#,16#0#,16#bc#,16#bc#,16#bc#,16#18#,16#18#,16#bc#,16#bc#,16#bc#,16#18#,16#14#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#9b#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#18#,16#bc#,16#18#,16#14#,16#bc#,16#bc#,16#bc#,16#18#,16#0#,16#bc#,16#bc#,16#bc#,16#18#,16#18#,16#bc#,16#bc#,16#bc#,16#18#,16#14#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#18#,16#bc#,16#14#,16#18#,16#bc#,16#bc#,16#b8#,16#18#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#20#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#0#,16#18#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#ff#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#ff#,16#ff#,16#bb#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#d7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#4#,16#fb#,16#20#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#ff#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#20#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#21#,16#d7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#1#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#4#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#0#,16#ff#,16#ff#,16#0#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#20#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#20#,16#0#,16#b7#,16#b7#,16#0#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#20#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#20#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#20#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#0#,16#4#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#4#,16#fb#,16#20#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#1#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#4#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#20#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#20#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#20#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#20#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#0#,16#d7#,16#d7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#0#,16#ff#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#0#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#ff#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#0#,16#ff#,16#ff#,16#9b#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#20#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#ff#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#9b#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#ff#,16#b7#,16#b7#,16#d7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#0#,16#18#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#0#,16#ff#,16#ff#,16#bb#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#9b#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#18#,16#18#,16#18#,16#18#,16#18#,16#14#,16#18#,16#18#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#b8#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#20#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#20#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#4#,16#fb#,16#20#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#9b#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#b8#,16#bc#,16#bc#,16#0#,16#18#,16#14#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#14#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#ff#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#d7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#bb#,16#ff#,16#0#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#0#,16#14#,16#18#,16#18#,16#14#,16#14#,16#18#,16#14#,16#18#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#b8#,16#bc#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#d7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#0#,16#18#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#1#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#14#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#0#,16#18#,16#18#,16#14#,16#14#,16#18#,16#18#,16#14#,16#18#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#4#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#0#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#14#,16#0#,16#18#,16#14#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#14#,16#18#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#20#,16#18#,16#14#,16#14#,16#14#,16#18#,16#18#,16#14#,16#14#,16#0#,16#14#,16#14#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#1#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#18#,16#18#,16#14#,16#18#,16#18#,16#18#,16#18#,16#14#,16#20#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#14#,16#18#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#4#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#0#,16#ff#,16#ff#,16#0#,16#ff#,16#4#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#14#,16#18#,16#14#,16#18#,16#14#,16#18#,16#18#,16#18#,16#0#,16#14#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#20#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#0#,16#b7#,16#b7#,16#0#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#0#,16#14#,16#18#,16#18#,16#18#,16#18#,16#18#,16#14#,16#18#,16#0#,16#18#,16#18#,16#18#,16#18#,16#14#,16#14#,16#18#,16#18#,16#18#,16#14#,16#18#,16#18#,16#18#,16#14#,16#14#,16#18#,16#18#,16#18#,16#18#,16#18#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#d7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#20#,16#18#,16#34#,16#18#,16#18#,16#18#,16#18#,16#18#,16#18#,16#0#,16#bc#,16#bc#,16#bc#,16#14#,16#14#,16#bc#,16#bc#,16#bc#,16#14#,16#18#,16#bc#,16#bc#,16#bc#,16#14#,16#14#,16#bc#,16#bc#,16#bc#,16#18#,16#18#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#18#,16#bc#,16#18#,16#18#,16#bc#,16#bc#,16#bc#,16#18#,16#0#,16#bc#,16#bc#,16#bc#,16#14#,16#14#,16#bc#,16#bc#,16#bc#,16#14#,16#18#,16#bc#,16#bc#,16#bc#,16#14#,16#14#,16#bc#,16#bc#,16#bc#,16#18#,16#18#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#0#,16#14#,16#bc#,16#18#,16#18#,16#bc#,16#bc#,16#b8#,16#14#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#0#,16#14#,16#bc#,16#bc#,16#bc#,16#bc#,16#b8#,16#bc#,16#bc#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#20#,16#0#,16#0#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#20#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#20#,16#bc#,16#bc#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#d7#,16#b7#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#20#,16#b8#,16#bc#,16#14#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#4#,16#fb#,16#20#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#20#,16#bc#,16#bc#,16#b8#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#bc#,16#bc#,16#bc#,16#b8#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#b8#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#1#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#bc#,16#bc#,16#18#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#4#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#20#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#b8#,16#bc#,16#bc#,16#bc#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#0#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#bc#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#d7#,16#0#,16#bc#,16#bc#,16#bc#,16#bc#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#20#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#bc#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d7#,16#b7#,16#b7#,16#0#,16#bc#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#0#,16#bc#,16#bc#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#0#,16#0#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#20#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#d7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#,16#d0#,16#fb#,16#fb#,16#fb#,16#fb#,16#fb#,16#0#,16#fb#,16#fb#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#fb#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#0#,16#d0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#fb#,16#fb#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#d7#,16#b7#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#,16#d0#,16#fb#,16#fb#,16#d0#,16#fb#,16#fb#,16#d0#,16#d0#,16#d0#,16#0#),
(16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#b7#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#,16#fb#,16#d0#,16#d0#,16#0#,16#d0#,16#d0#,16#d0#,16#d0#,16#d0#,16#0#));