type memoryPicture is array(0 to 30, 0 to 14) of integer;
constant picture : memoryPicture:=(
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#0#,16#0#,16#ff#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#0#,16#0#,16#ff#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#ff#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#ff#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#ff#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#ff#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#0#,16#0#,16#ff#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#0#,16#0#,16#ff#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#));