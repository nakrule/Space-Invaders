type memoryPicture is array(0 to 179, 0 to 108) of integer;
constant picture : memoryPicture:=(
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#92#,16#b6#,16#db#,16#ff#,16#ff#,16#ff#,16#db#,16#db#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#24#,16#92#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#24#,16#0#,16#6e#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6e#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#25#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#49#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#49#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#24#,16#0#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#49#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#49#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#92#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#92#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#49#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#49#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#25#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#92#,16#0#,16#0#,16#0#,16#92#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6e#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#25#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#92#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#6d#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6d#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6e#,16#49#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#6d#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6e#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#24#,16#49#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#25#,16#0#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#24#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#0#,16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#25#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6e#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#db#,16#b6#,16#92#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#),
(16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6d#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#),
(16#0#,16#0#,16#0#,16#0#,16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#49#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#0#,16#0#,16#24#,16#b6#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#24#,16#0#,16#24#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#25#,16#49#,16#92#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#b6#,16#92#,16#92#,16#92#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#49#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#24#,16#0#,16#25#,16#0#,16#24#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#49#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6e#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6e#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#25#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#49#,16#24#,16#0#,16#0#,16#25#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#49#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#6e#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#6d#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#6d#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#49#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#24#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#0#,16#0#,16#49#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#6e#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#92#,16#0#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#25#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#24#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#49#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6d#,16#0#,16#0#,16#0#,16#25#,16#0#,16#25#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#0#,16#0#,16#0#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#24#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#da#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6d#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6e#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#24#,16#0#,16#24#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#da#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#25#,16#24#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#24#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#24#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#24#,16#0#,16#24#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#0#),
(16#0#,16#0#,16#0#,16#49#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#24#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#25#,16#0#,16#24#,16#0#,16#24#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#0#,16#25#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#49#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#b6#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#6d#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#24#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#49#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#92#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#25#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#24#,16#92#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#24#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#92#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#24#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#24#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#92#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#25#,16#0#,16#0#,16#24#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6e#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#0#,16#0#,16#24#,16#6e#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#92#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6e#,16#24#,16#24#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#24#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#25#,16#24#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6d#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#6d#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#6e#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6d#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#24#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#6d#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6e#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#24#,16#24#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#6d#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#24#,16#49#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6e#,16#0#,16#25#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#24#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#92#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#24#,16#24#,16#0#,16#0#,16#92#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#25#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#24#,16#0#,16#92#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#24#,16#24#,16#0#,16#0#,16#6d#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#92#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#6d#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#6d#,16#0#,16#25#,16#25#,16#0#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#24#,16#b6#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#6e#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#49#,16#0#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#25#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#25#,16#24#,16#0#,16#24#,16#0#,16#0#,16#25#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#25#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#92#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#92#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#49#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#49#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#b6#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#49#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#24#,16#24#,16#0#,16#49#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#24#,16#0#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#25#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#24#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#49#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#24#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#24#,16#0#,16#24#,16#49#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#b6#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#25#,16#db#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#92#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#24#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#24#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#92#,16#ff#,16#ff#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#25#,16#0#,16#24#,16#0#),
(16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#ff#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#));