----------------------------------------------------------------------------------
-- Company:        HES-SO
-- Engineer:       Samuel Riedo & Pascal Roulin
-- Create Date:    11:24:52 03/02/2017
-- Design Name:    SpaceInvadersPackage.vhd
-- Project Name:   Space Invaders - FPGA Edition
-- Target Devices: Digilent NEXYS 3 (Xilinx Spartan 6 XC6LX16-CS324)
-- Description:    Contain all constant.
-- Revision 0.01 - File Created
--          1.00 - Add VGA contants
--          1.1  - Add Inputs contants
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package SpaceInvadersPackage is

----------------------------------------------------------------------------------
  -- VGA
  constant HMAX             : integer := 1056;
  constant VMAX             : integer := 628;
  constant HLINES           : integer := 800;
  constant VLINES           : integer := 600;
  constant HSP              : integer := 968;
  constant HFP              : integer := 840;
  constant VFP              : integer := 601;
  constant VSP              : integer := 605;
  ----------------------------------------------------------------------------------
  -- Inputs
  constant fireSpeed        : integer := 600000;
  constant shipSpeed        : integer := 100000;
  constant alienSpeed       : integer := 6000000;
  constant maxShipPosValue  : integer := 736;  -- must be pair
  constant shipMargin       : integer := 50;   -- minimum space between side screen and ship
  constant alienXMargin     : integer := 50;   -- minimum space between side screen and aliens
  constant alienYUpMargin   : integer := 50;   -- minimum space between top screen and aliens
  constant alienYDownMargin : integer := 200;  -- maximum space between top screen and aliens
  constant maxAlienJump     : integer := 10;   -- max pixel aliens can shift in a single time
----------------------------------------------------------------------------------
  -- rocketManager
	constant missileSpeed    : integer := 60000; -- missile speed
	constant rocketLength	 : integer := 10;    -- rocket length in pixel
	constant rocketColor     : std_logic_vector(7 downto 0) := "11111111";
----------------------------------------------------------------------------------
  -- Tables of aliens and ship

  -- 0 = no alien
  -- 1 = blue, 3 = dark blue, 5 = green, 7 = purple, 9 = yellow
  -- 2 = blue alien killed, 4 = dark blue alien killed, etc ...
  type aliensArray is array(9 downto 0, 4 downto 0) of integer range 0 to 10;
  signal aliens : aliensArray := (others => (others => 1));  -- Initialized to 0

  -- All aliens are 30x30
  type alienPicture is array(0 to 29, 0 to 29) of integer;

  constant blueAlien : alienPicture := (
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#21#, 16#21#, 16#4#, 16#4#, 16#4#, 16#4#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#21#, 16#21#, 16#4#, 16#4#, 16#4#, 16#4#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#21#, 16#21#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#21#, 16#21#, 16#0#, 16#0#),
    (16#20#, 16#20#, 16#4#, 16#4#, 16#0#, 16#0#, 16#24#, 16#24#, 16#56#, 16#56#, 16#77#, 16#77#, 16#56#, 16#56#, 16#76#, 16#76#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#1#, 16#20#, 16#20#),
    (16#20#, 16#20#, 16#4#, 16#4#, 16#0#, 16#0#, 16#24#, 16#24#, 16#56#, 16#56#, 16#77#, 16#77#, 16#56#, 16#56#, 16#76#, 16#76#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#5#, 16#4#, 16#0#, 16#0#, 16#20#, 16#20#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#1#, 16#1#, 16#21#, 16#21#, 16#0#, 16#0#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#0#, 16#0#, 16#76#, 16#76#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#1#, 16#1#, 16#21#, 16#21#, 16#0#, 16#0#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#0#, 16#0#, 16#76#, 16#76#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#21#, 16#21#, 16#24#, 16#24#, 16#76#, 16#76#, 16#0#, 16#20#, 16#76#, 16#76#, 16#77#, 16#77#, 16#56#, 16#56#, 16#76#, 16#76#, 16#76#, 16#76#, 16#20#, 16#20#, 16#0#, 16#1#, 16#21#, 16#21#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#21#, 16#21#, 16#24#, 16#24#, 16#76#, 16#76#, 16#0#, 16#0#, 16#76#, 16#76#, 16#77#, 16#77#, 16#56#, 16#56#, 16#76#, 16#76#, 16#76#, 16#76#, 16#20#, 16#20#, 16#0#, 16#0#, 16#21#, 16#21#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#76#, 16#76#, 16#76#, 16#76#, 16#0#, 16#0#, 16#76#, 16#76#, 16#76#, 16#76#, 16#0#, 16#0#, 16#0#, 16#0#, 16#4#, 16#1#, 16#0#, 16#0#, 16#0#, 16#0#, 16#4#, 16#4#),
    (16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#76#, 16#76#, 16#76#, 16#76#, 16#0#, 16#0#, 16#76#, 16#76#, 16#76#, 16#76#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#4#, 16#4#),
    (16#0#, 16#0#, 16#24#, 16#24#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#77#, 16#77#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#24#, 16#24#, 16#20#, 16#20#, 16#1#, 16#1#),
    (16#0#, 16#0#, 16#24#, 16#24#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#77#, 16#77#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#24#, 16#24#, 16#20#, 16#20#, 16#0#, 16#1#),
    (16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#20#, 16#20#, 16#0#, 16#1#, 16#0#, 16#0#, 16#4#, 16#0#, 16#0#, 16#0#, 16#1#, 16#1#),
    (16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#1#, 16#1#),
    (16#20#, 16#20#, 16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#77#, 16#77#, 16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#21#, 16#21#),
    (16#20#, 16#20#, 16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#77#, 16#77#, 16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#21#),
    (16#0#, 16#1#, 16#20#, 16#20#, 16#0#, 16#0#, 16#20#, 16#20#, 16#56#, 16#56#, 16#76#, 16#76#, 16#21#, 16#1#, 16#76#, 16#76#, 16#76#, 16#76#, 16#4#, 16#4#, 16#20#, 16#20#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#20#, 16#20#, 16#56#, 16#56#, 16#76#, 16#76#, 16#1#, 16#1#, 16#76#, 16#76#, 16#76#, 16#76#, 16#4#, 16#4#, 16#20#, 16#20#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#1#, 16#0#, 16#76#, 16#76#, 16#4#, 16#4#, 16#76#, 16#76#, 16#56#, 16#56#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#76#, 16#76#, 16#4#, 16#4#, 16#76#, 16#76#, 16#56#, 16#56#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#),
    (16#4#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#20#, 16#20#, 16#76#, 16#76#, 16#77#, 16#77#, 16#77#, 16#77#, 16#0#, 16#0#, 16#77#, 16#76#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#4#, 16#4#, 16#20#, 16#20#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#20#, 16#20#, 16#76#, 16#76#, 16#77#, 16#77#, 16#77#, 16#77#, 16#0#, 16#0#, 16#77#, 16#76#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#1#, 16#0#, 16#0#, 16#0#, 16#0#, 16#4#, 16#20#, 16#20#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#4#, 16#20#, 16#20#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#4#, 16#4#, 16#20#, 16#20#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#76#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#21#, 16#21#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#1#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#21#, 16#21#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#1#, 16#1#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#1#, 16#1#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#1#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#));

  constant darkBlueAlien : alienPicture := (
    (16#0#, 16#0#, 16#0#, 16#0#, 16#1#, 16#1#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#1#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#1#, 16#1#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#20#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#4#, 16#24#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#));

  constant greenAlien : alienPicture := (
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#98#, 16#98#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#98#, 16#98#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#98#, 16#98#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#98#, 16#98#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#98#, 16#98#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#98#, 16#98#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#98#, 16#98#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#98#, 16#98#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#98#, 16#98#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#98#, 16#98#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#98#, 16#98#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#98#, 16#98#, 16#98#, 16#98#, 16#0#, 16#0#, 16#98#, 16#98#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#));

  constant purpleAlien : alienPicture := (
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#21#, 16#21#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#21#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c7#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#c3#, 16#c3#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#21#, 16#21#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#21#, 16#21#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#));

  constant yellowAlien : alienPicture := (
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#1#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#4#, 16#4#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#20#, 16#20#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#fc#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#20#, 16#20#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#));


  type shipPicture is array(0 to 61, 0 to 29) of integer;
  constant ship : shipPicture := (
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#),
    (16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#, 16#0#));
----------------------------------------------------------------------------------
end SpaceInvadersPackage;
