type memoryPicture is array(0 to 29, 0 to 29) of integer;
constant picture : memoryPicture:=(
(16#0#,16#0#,16#0#,16#0#,16#1#,16#1#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#1#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#1#,16#1#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#4#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#4#,16#4#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#20#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#20#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#3#,16#3#,16#3#,16#3#,16#3#,16#3#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#20#,16#20#,16#20#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#20#,16#20#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#),
(16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#4#,16#24#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#,16#0#));